//**********************************************************************
//  Project: ASIC-Hw4
//  File: half_adder.v
//  Description: half adder
//  Author: Ruiqi Tang
//  Timestamp:
//----------------------------------------------------------------------
// Code Revision History:
// Ver:     | Author    | Mod. Date     | Changes Made:
// v1.0.0   | R.T.      | 2024/04/18    | Initial version
//**********************************************************************


module half_adder(
    a,
    enable,
    sum,
    c_out
);

//**********************************************************************
// --- Parameter
//**********************************************************************
    parameter DATAWIDTH = 8;

//**********************************************************************
// --- Input/Output Declaration
//**********************************************************************
    input  wire  [DATAWIDTH-1:0]    a;
    input  wire                     enable;
    output wire  [DATAWIDTH-1:0]    sum;
    output wire                     c_out;

//**********************************************************************
// --- Main Core
//**********************************************************************
    assign {c_out, sum} = enable ? (a + 1'b1) : ({1'b0, {(DATAWIDTH-1){1'bz}}});

endmodule